
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_std.all;
use work.SADlibrary.all;


entity testbench is

end testbench;


architecture tb of testbench is

    constant data_width                                 : integer := 16;
    constant matrix_size                                : std_logic_vector(data_width - 1 downto 0) := x"0010";
    signal clk, rst, start, w_en_x, w_en_y, done        : std_logic;
    signal x_in, y_in, SAD_o                            : std_logic_vector(data_width - 1 downto 0);

    begin
        computeSAD_process  : computeSAD  generic map(data_width, matrix_size)
                                             port map(clk, rst, start, w_en_x, w_en_y, x_in, y_in, SAD_o, done);

        clock_sig:
            process 
                begin  
                    clk <= '0';
                    wait for 1 ns;
                    clk <= '1';
                    wait for 1 ns;
            end process;
        


        reset:
            process
                begin
                    rst <= '1';
                    wait for 4 ns;
                    rst <= '0';
                    wait;
            end process;
        
        write_enable_x:
            process 
                begin 
                    w_en_x <= '0';
                    wait for 5 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 400 ns;
                    w_en_x <= '0';
                    wait for 5 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait for 2 ns;
                    w_en_x <= '1';
                    wait for 2 ns;
                    w_en_x <= '0';
                    wait;
            end process;

        write_enable_y:
            process 
                begin 
                    w_en_y <= '0';
                    wait for 5 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    --wait for 2 ns;
                    wait for 400 ns;
                    w_en_y <= '0';
                    wait for 5 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait for 2 ns;
                    w_en_y <= '1';
                    wait for 2 ns;
                    w_en_y <= '0';
                    wait;
            end process;
        
        compute:
            process
                begin
                    start <= '0';
                    wait for 5 ns;
                    x_in <= x"F4F3";
                    y_in <= x"0001";
                    wait for 4 ns;
                    x_in <= x"0012";
                    y_in <= x"000B";
                    wait for 4 ns;
                    x_in <= x"0009";
                    y_in <= x"0001";
                    wait for 4 ns;
                    x_in <= x"FF2F";
                    y_in <= x"000A";
                    wait for 4 ns;
                    x_in <= x"0007";
                    y_in <= x"FFFF";
                    wait for 4 ns;
                    x_in <= x"0B02";
                    y_in <= x"0012";
                    wait for 4 ns;
                    x_in <= x"0002";
                    y_in <= x"0006";
                    wait for 4 ns;
                    x_in <= x"00F6";
                    y_in <= x"000B";
                    wait for 4 ns;
                    x_in <= x"0C05";
                    y_in <= x"0001";
                    wait for 4 ns;
                    x_in <= x"FFFA";
                    y_in <= x"00DD";
                    wait for 4 ns;
                    x_in <= x"000C";
                    y_in <= x"00BB";
                    wait for 4 ns;
                    x_in <= x"000A";
                    y_in <= x"0A09";
                    wait for 4 ns;
                    x_in <= x"00D8";
                    y_in <= x"0000";
                    wait for 4 ns;
                    x_in <= x"000F";
                    y_in <= x"000F";
                    wait for 4 ns;
                    x_in <= x"0012";
                    y_in <= x"FFF7";
                    wait for 4 ns;
                    x_in <= x"FFFF";
                    y_in <= x"0000";
                    wait for 2 ns;
                    start <= '1';
                    wait for 400 ns;
                    start <= '0';
                    wait for 5 ns;
                    -- TEST 2
                    x_in <= x"FFF3";
                    y_in <= x"00AA";
                    wait for 4 ns;
                    x_in <= x"0010";
                    y_in <= x"00DB";
                    wait for 4 ns;
                    x_in <= x"00DD";
                    y_in <= x"FFA9";
                    wait for 4 ns;
                    x_in <= x"0069";
                    y_in <= x"0021";
                    wait for 4 ns;
                    x_in <= x"00E7";
                    y_in <= x"FF11";
                    wait for 4 ns;
                    x_in <= x"0B0E";
                    y_in <= x"0112";
                    wait for 4 ns;
                    x_in <= x"0102";
                    y_in <= x"000A";
                    wait for 4 ns;
                    x_in <= x"FFF6";
                    y_in <= x"000B";
                    wait for 4 ns;
                    x_in <= x"FFF5";
                    y_in <= x"FFB1";
                    wait for 4 ns;
                    x_in <= x"FFFA";
                    y_in <= x"FFDD";
                    wait for 4 ns;
                    x_in <= x"FF1C";
                    y_in <= x"FFFB";
                    wait for 4 ns;
                    x_in <= x"000A";
                    y_in <= x"0A09";
                    wait for 4 ns;
                    x_in <= x"00D8";
                    y_in <= x"FEE0";
                    wait for 4 ns;
                    x_in <= x"FFEF";
                    y_in <= x"0020";
                    wait for 4 ns;
                    x_in <= x"0A12";
                    y_in <= x"0007";
                    wait for 4 ns;
                    x_in <= x"FFF0";
                    y_in <= x"000C";
                    wait for 2 ns;
                    start <= '1';
                    wait;

            end process;


end tb;